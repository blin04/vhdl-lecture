library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package constants is
    constant CLK_PERIOD : time := 50 ns;
end package;
